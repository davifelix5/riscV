module program_counter (
    // Sinais de controle
    input CLK,
    input LOAD,
    input RST,
    input wire pc_next_sel,
    input wire pc_adder_sel,
    // Valores da instrução
    input wire[63:0] immediate,
    input wire[6:0] opcode,
    input wire[2:0] func,
    // Saída do regfile
    input wire[63:0] Dout_rs1,
    // Flags
    input wire EQ,
    input wire LT_SN,
    input wire LT_UN,
    input wire GT_SN,
    input wire GT_UN,
    // Endereço da memória de instruções
    output wire [63:0] addr,
    output wire[63:0] pc_to_store
);

    reg sel;

    always @(*) begin
        case (func)
            3'b000: sel = EQ;
            3'b001: sel = ~EQ;
            3'b100: sel = LT_SN;
            3'b101: sel = GT_SN;
            3'b110: sel = LT_UN;
            3'b111: sel = GT_UN;
            default: sel = 0;
        endcase
    end

    wire[63:0] pc_next, pc_adder, primary_adder_res, secondary_adder_res;
    wire final_pc_adder_sel, final_pc_next_sel;

    // Para que sel seja utilizado, opcode tem que ser 1100011
    assign final_pc_next_sel = opcode == 7'b1100011 ? sel : pc_next_sel;
    assign final_pc_adder_sel = opcode == 7'b1100011 ? 1'b1 : pc_adder_sel; 

    assign pc_adder = final_pc_adder_sel ? addr : Dout_rs1;
    assign pc_next = final_pc_next_sel ? secondary_adder_res : primary_adder_res;
    assign pc_to_store = primary_adder_res;
    

    adder #(.SIZE(64)) primary_adder (
        .X(addr),
        .Y(64'd4),
        .Cin(1'b0),
        .S(primary_adder_res)
    );

    adder #(.SIZE(64)) secondary_adder (
        .X(immediate),
        .Y(pc_adder),
        .Cin(1'b0),
        .S(secondary_adder_res)
    );

    register_negedge_with_reset #(.SIZE(64)) PC (.IN(pc_next), .OUT(addr), .RST(RST), .LOAD(LOAD), .CLK(CLK));

endmodule